`timescale 1ns / 1ps

module ROM (
    input  logic [31:0] addr,
    output logic [31:0] data
);
    logic [31:0] rom[0:2**8-1];

    initial begin
        $readmemh("code.mem", rom);

//========================================STORE=================================================
        // rom[0]  = 32'h04002023; // sw   x0,  0x40(x0)   ; mem[0x40..0x43]=0
        // rom[1]  = 32'h04002223; // sw   x0,  0x44(x0)   ; mem[0x44..0x47]=0
        // rom[2]  = 32'h04002423; // sw   x0,  0x48(x0)   ; mem[0x48..0x4B]=0

        // //  SB 검증: 각 바이트 lane에 0x11,22,33,44
        // rom[3]  = 32'h01100513; // addi x10, x0, 0x11
        // rom[4]  = 32'h02200593; // addi x11, x0, 0x22
        // rom[5]  = 32'h03300613; // addi x12, x0, 0x33
        // rom[6]  = 32'h04400693; // addi x13, x0, 0x44
        // rom[7]  = 32'h04a00023; // sb   x10, 0x40(x0)   ; lane0 -> [0x40]=11
        // rom[8]  = 32'h04b000a3; // sb   x11, 0x41(x0)   ; lane1 -> [0x41]=22
        // rom[9]  = 32'h04c00123; // sb   x12, 0x42(x0)   ; lane2 -> [0x42]=33
        // rom[10] = 32'h04d001a3; // sb   x13, 0x43(x0)   ; lane3 -> [0x43]=44
        // rom[11] = 32'h04002a03; // lw   x20,0x40(x0)    ; x20=0x44332211 (검증)

        // //  SH 검증: 하위=0x5566, 상위=0x7788
        // rom[12] = 32'h00005737; // lui  x14, 0x00005
        // rom[13] = 32'h56670713; // addi x14, x14, 0x566 ; x14=0x00005566
        // rom[14] = 32'h000077b7; // lui  x15, 0x00007
        // rom[15] = 32'h78878793; // addi x15, x15, 0x788 ; x15=0x00007788

        // rom[16] = 32'h04002223; // sw   x0,  0x44(x0)   ; 다시 0으로
        // rom[17] = 32'h04e01223; // sh   x14, 0x44(x0)   ; 하위 하프 0x5566
        // rom[18] = 32'h04f01323; // sh   x15, 0x46(x0)   ; 상위 하프 0x7788
        // rom[19] = 32'h04402a83; // lw   x21,0x44(x0)    ; x21=0x77885566 (검증)

        // //  SW 검증: 0xA1B2C3D4
        // rom[20] = 32'ha1b2c837; // lui  x16, 0xA1B2C
        // rom[21] = 32'h3d480813; // addi x16, x16, 0x3D4 ; x16=0xA1B2C3D4
        // rom[22] = 32'h05002423; // sw   x16, 0x48(x0)
        // rom[23] = 32'h04802b03; // lw   x22, 0x48(x0)   ; x22=0xA1B2C3D4 (검증)

//========================================Load=================================================

        // // 0으로 초기화
        // rom[0]  = 32'h04002023; // sw x0, 0x40(x0)  ; [0x40..43]=0
        // rom[1]  = 32'h04002223; // sw x0, 0x44(x0)  ; [0x44..47]=0
        // rom[2]  = 32'h04002423; // sw x0, 0x48(x0)  ; [0x48..4B]=0
        
        // //  LB용 바이트 : [0x40]=7F, [0x41]=80, [0x42]=01, [0x43]=F2
        // rom[3]  = 32'h07F00513; // addi x10,x0,0x7F
        // rom[4]  = 32'h08000593; // addi x11,x0,0x80
        // rom[5]  = 32'h00100613; // addi x12,x0,0x01
        // rom[6]  = 32'h0F200693; // addi x13,x0,0xF2
        // rom[7]  = 32'h04A00023; // sb   x10,0x40(x0)  ; lane0
        // rom[8]  = 32'h04B000A3; // sb   x11,0x41(x0)  ; lane1
        // rom[9]  = 32'h04C00123; // sb   x12,0x42(x0)  ; lane2
        // rom[10] = 32'h04D001A3; // sb   x13,0x43(x0)  ; lane3
        
        // //  LB 4케이스 로드(부호확장 확인)
        // rom[11] = 32'h04000A03; // lb x20,0x40(x0)  ; x20=0x0000007F
        // rom[12] = 32'h04100A83; // lb x21,0x41(x0)  ; x21=0xFFFFFF80
        // rom[13] = 32'h04200B03; // lb x22,0x42(x0)  ; x22=0x00000001
        // rom[14] = 32'h04300B83; // lb x23,0x43(x0)  ; x23=0xFFFFFFF2
        
        // // ── LH용 하프워드 : 하위=0x7F7F(양수), 상위=0x8001(음수)
        // rom[15] = 32'h00008737; // lui  x14,0x00008      ; x14=0x00008000
        // rom[16] = 32'hF7F70713; // addi x14,x14,-129     ; x14=0x00007F7F
        // rom[17] = 32'h000087B7; // lui  x15,0x00008      ; x15=0x00008000
        // rom[18] = 32'h00178793; // addi x15,x15,1        ; x15=0x00008001
        // rom[19] = 32'h04E01223; // sh   x14,0x44(x0)     ; [0x44..45]=7F 7F
        // rom[20] = 32'h04F01323; // sh   x15,0x46(x0)     ; [0x46..47]=01 80
        
        // //  LH 2케이스 로드(부호확장 확인)
        // rom[21] = 32'h04401C03; // lh x24,0x44(x0)  ; x24=0x00007F7F
        // rom[22] = 32'h04601C83; // lh x25,0x46(x0)  ; x25=0xFFFF8001
        
        // //  LW용 워드 
        // rom[23] = 32'hA1B2C837; // lui  x16,0xA1B2C      ; x16=0xA1B2C000
        // rom[24] = 32'h3D480813; // addi x16,x16,0x3D4    ; x16=0xA1B2C3D4
        // rom[25] = 32'h05002423; // sw   x16,0x48(x0)     ; 
        
        // //  LW 로드 
        // rom[26] = 32'h04802D03; // lw  x26,0x48(x0) ; x26=0xA1B2C3D4

        // //  LBU 4케이스 (제로확장 확인): [0x40]=7F, [0x41]=80, [0x42]=01, [0x43]=F2
        // rom[27] = 32'h04004B83; // lbu x23,0x40(x0) ; 기대: x23=0x0000007F
        // rom[28] = 32'h04104C03; // lbu x24,0x41(x0) ; 기대: x24=0x00000080
        // rom[29] = 32'h04204C83; // lbu x25,0x42(x0) ; 기대: x25=0x00000001
        // rom[30] = 32'h04304D03; // lbu x26,0x43(x0) ; 기대: x26=0x000000F2

        // //  LHU 2케이스 (제로확장 확인)
        // rom[31] = 32'h04405D83; // lhu x27,0x44(x0) ; 기대: x27=0x00007F7F
        // rom[32] = 32'h04605E03; // lhu x28,0x46(x0) ; 기대: x28=0x00008001

//==============================================Branch=========================================
  
    // //  BEQ: x2를 0→1→2로 만들며, x2==x1(=1)일 때만 1번 루프 
    // rom[0]  = 32'h00100093; // addi x1, x0, 1
    // rom[1]  = 32'h00000113; // addi x2, x0, 0
    // rom[2]  = 32'h00110113; // L_BEQ: addi x2, x2, 1
    // rom[3]  = 32'hfe110ee3; // beq  x2, x1, L_BEQ   ; offset -4
    
    // //  BNE: x3를 0→1→2, x4=2. x3!=x4일 때만 루프(1회) 
    // rom[4]  = 32'h00200213; // addi x4, x0, 2
    // rom[5]  = 32'h00000193; // addi x3, x0, 0
    // rom[6]  = 32'h00118193; // L_BNE: addi x3, x3, 1
    // rom[7]  = 32'hfe419ee3; // bne  x3, x4, L_BNE   ; -4
    
    // //  BLT(signed): x5를 0→1→2, x6=2. x5<x6일 때 루프(1회) 
    // rom[8]  = 32'h00200313; // addi x6, x0, 2
    // rom[9]  = 32'h00000293; // addi x5, x0, 0
    // rom[10] = 32'h00128293; // L_BLT: addi x5, x5, 1
    // rom[11] = 32'hfe62cee3; // blt  x5, x6, L_BLT   ; -4
    
    // //  BGE(signed): x7=2부터 1→0→-1, x7>=0일 때 루프(2회) 
    // rom[12] = 32'h00200393; // addi x7, x0, 2
    // rom[13] = 32'hfff38393; // L_BGE: addi x7, x7, -1
    // rom[14] = 32'hfe03dee3; // bge  x7, x0, L_BGE   ; -4
    
    // //  BLTU(unsigned): x8 0→1→2, x9=2. x8<x9일 때 루프(1회) 
    // rom[15] = 32'hFFE00493; // addi x9, x0, -2
    // rom[16] = 32'h00000413; // addi x8, x0, 0
    // rom[17] = 32'h00140413; // L_BLTU: addi x8, x8, 1
    // rom[18] = 32'hfe946ee3; // bltu x8, x9, L_BLTU  ; -4
    
    // //  BGEU(unsigned): x10=2부터 1→0, x11=1. x10>=x11일 때 루프(1회) 
    // rom[19] = 32'h00100593; // addi x11, x0, 1
    // rom[20] = 32'h00200513; // addi x10, x0, 2
    // rom[21] = 32'hfff50513; // L_BGEU: addi x10, x10, -1
    // rom[22] = 32'hfeb57ee3; // bgeu x10, x11, L_BGEU ; -4

//==========================================================================================
        // // R-Type  funct7(7) | rs2(5) | rs1(5) | funct3(3) | rd(5) | opcode(7)
        // rom[0] = 32'b0000000_00001_00010_000_00100_0110011;  // add  x4,  x2, x1         
        // rom[1] = 32'b0100000_00001_00010_000_00101_0110011;  // sub  x5,  x2, x1
        // rom[2] = 32'b0000000_00001_00010_001_00110_0110011;  // sll  x6,  x2, x1
        // rom[3] = 32'b0000000_00001_00010_101_00111_0110011;  // srl  x7,  x2, x1
        // rom[4] = 32'b0100000_00001_00010_101_01000_0110011;  // sra  x8,  x2, x1
        // rom[5] = 32'b0000000_00001_00010_010_01001_0110011;  // slt  x9,  x2, x1
        // rom[6] = 32'b0000000_00001_00010_011_01010_0110011;  // sltu x10, x2, x1
        // rom[7] = 32'b0000000_00001_00010_100_01011_0110011;  // xor  x11, x2, x1
        // rom[8] = 32'b0000000_00001_00010_110_01100_0110011;  // or   x12, x2, x1
        // rom[9] = 32'b0000000_00001_00010_111_01101_0110011;  // and  x13, x2, x1    
        
        // // S-Type  imm[11:5](7) | rs2(5) | rs1(5) | funct3(3) | imm[4:0](5) | opcode(7)  
        // rom[10] = 32'b0000000_00100_00000_010_10000_0100011; // sw x4, 16(x0)         
        // rom[11] = 32'b0000000_00100_00000_000_10100_0100011; // sb x4, 20(x0)
        // rom[12] = 32'b0000000_00100_00000_001_11000_0100011; // sh x4, 24(x0)    

        // // L-Type  imm[11:0](12) | rs1(5) | funct3(3) | rd(5) | opcode(7)
        // rom[13] = 32'b000000010000_00000_010_01110_0000011;  // lw  x14, 16(x0)
        // rom[14] = 32'b000000010100_00000_000_01111_0000011;  // lb  x15, 20(x0)        
        // rom[15] = 32'b000000011000_00000_001_10000_0000011;  // lh  x16, 24(x0)
        // rom[16] = 32'b000000010100_00000_100_10001_0000011;  // lbu x17, 20(x0)
        // rom[17] = 32'b000000011000_00000_101_10010_0000011;  // lhu x18, 24(x0)

        // // I-Type  imm[11:0](12) | rs1(5) | funct3(3) | rd(5) | opcode(7)
        // rom[18] = 32'b111111111000_00010_000_10011_0010011;  // addi  x19, x2, -8       
        // rom[19] = 32'b111111111100_00010_010_10100_0010011;  // slti  x20, x2, -4
        // rom[20] = 32'b111111111100_00010_011_10101_0010011;  // sltiu x21, x2, -4
        // rom[21] = 32'b000000000100_00010_100_10110_0010011;  // xori  x22, x2,  4 
        // rom[22] = 32'b000000000100_00010_110_10111_0010011;  // ori   x23, x2,  4 
        // rom[23] = 32'b000000000100_00010_111_11000_0010011;  // andi  x24, x2,  4 
        // rom[24] = 32'b0000000_00001_00010_001_11001_0010011; // slli  x25, x2,  1
        // rom[25] = 32'b0000000_00001_00100_101_11010_0010011; // srli  x26, x4,  1
        // rom[26] = 32'b0100000_00001_00100_101_11011_0010011; // srai  x27, x4,  1

        // // B-Type  imm[12|10:5](7) | rs2(5) | rs1(5) | funct3(3) | imm[4:1|114(5) | opcode(7)
        // rom[27] = 32'b0000000_00010_00011_000_00100_1100011; // beq  x3, x2, 4
        // rom[28] = 32'b0000000_00010_00011_001_00100_1100011; // bne  x3, x2, 4
        // rom[29] = 32'b0000000_00010_00011_100_00100_1100011; // blt  x3, x2, 4 
        // rom[30] = 32'b0000000_00010_00011_101_00100_1100011; // bge  x3, x2, 4 
        // rom[31] = 32'b0000000_00010_00011_110_00100_1100011; // bltu x3, x2, 4 
        // rom[32] = 32'b0000000_00010_00011_111_00100_1100011; // bgeu x3, x2, 4     

        // // U-Type  imm[31:12](20) | rd(5) | opcode(7)
        // rom[33] = 32'b00000000000000000001_11100_0110111;    // lui x28, 1          
        // rom[34] = 32'b00000000000000000001_11101_0010111;    // auipc x29, 1

        // // J-Type  imm[20|10:1|11|19:12](20) | rd(5) | opcode(7)
        // rom[35] = 32'b0_0000000010_0_00000000_11110_1101111; // jal x30, 4

        // // J-Type (JALR)  imm[11:0](12) | rs1(5) | funct3(3) | rd(5) | opcode(7)
        // rom[36] = 32'b000000000100_00100_000_11111_1100111;  // jalr x31, x4, 4
    
    end

    assign data = rom[addr[31:2]];
endmodule


